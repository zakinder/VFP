-------------------------------------------------------------------------------
--
-- Filename    : recolor_space_cluster.vhd
-- Create Date : 05062019 [05-06-2019]
-- Author      : Zakinder
--
-- Description:
-- This file instantiation
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.fixed_pkg.all;
use work.float_pkg.all;
use work.constants_package.all;
use work.vpf_records.all;
use work.vfp_pkg.all;
use work.ports_package.all;
entity recolor_space_cluster is
generic (
    neighboring_pixel_threshold : integer := 255;
    img_width                   : integer := 1920;
    i_data_width                : integer := 8);
port (
    clk                         : in  std_logic;
    reset                       : in  std_logic;
    iRgb                        : in channel;
    txCord                      : in coord;
    oRgb                        : out channel);
end recolor_space_cluster;
architecture behavioral of recolor_space_cluster is
    signal re_00_space     : channel;
    signal re_01_space     : channel;
    signal re_02_space     : channel;
    signal re_03_space     : channel;
    signal re_04_space     : channel;
    signal re_05_space     : channel;
    signal re_06_space     : channel;
    signal re_07_space     : channel;
    signal re_08_space     : channel;
    signal re_09_space     : channel;
    signal re_10_space     : channel;
    signal re_11_space     : channel;
    signal re_12_space     : channel;
    signal re_13_space     : channel;
    signal re_14_space     : channel;
    signal re_15_space     : channel;
    signal re_16_space     : channel;
    signal re_17_space     : channel;
    signal re_18_space     : channel;
    signal re_19_space     : channel;
    signal re_20_space     : channel;
    signal re_21_space     : channel;
    signal re_22_space     : channel;
    signal re_23_space     : channel;
    signal re_24_space     : channel;
begin 
------------------------------------------------------------------------------
recolor_space_1_inst: pixel_localization
generic map(
    neighboring_pixel_threshold => 10,
    img_width                   => img_width,
    i_data_width                => i_data_width)
port map(
    clk                => clk,
    reset              => reset,
    iRgb               => iRgb,
    txCord             => txCord,
    oRgb               => re_00_space);
rgb_contrast_brightness_1_inst: rgb_contrast_brightness_level_1
generic map (
    contrast_val  => to_sfixed(0.90,16,-3),
    exposer_val  => 0)
port map (                  
    clk               => clk,
    rst_l             => reset,
    iRgb              => re_00_space,
    oRgb              => re_01_space);
rgb_range_1_inst: rgb_range
generic map (
    i_data_width       => i_data_width)
port map (                  
    clk                => clk,
    reset              => reset,
    iRgb               => re_01_space,
    oRgb               => re_02_space);
------------------------------------------------------------------------------
------------------------------------------------------------------------------
recolor_space_2_inst: pixel_localization
generic map(
    neighboring_pixel_threshold => 12,
    img_width                   => img_width,
    i_data_width                => i_data_width)
port map(
    clk                => clk,
    reset              => reset,
    txCord             => txCord,
    iRgb               => re_02_space,
    oRgb               => re_03_space);
rgb_contrast_brightness_2_inst: rgb_contrast_brightness_level_1
generic map (
    contrast_val  => to_sfixed(1.20,16,-3),
    exposer_val  => 0)
port map (                  
    clk               => clk,
    rst_l             => reset,
    iRgb              => re_03_space,
    oRgb              => re_04_space);
rgb_range_2_inst: rgb_range
generic map (
    i_data_width       => i_data_width)
port map (                  
    clk                => clk,
    reset              => reset,
    iRgb               => re_04_space,
    oRgb               => re_05_space);
------------------------------------------------------------------------------
------------------------------------------------------------------------------
recolor_space_3_inst: pixel_localization
generic map(
    neighboring_pixel_threshold => 13,
    img_width         => img_width,
    i_data_width      => i_data_width)
port map(
    clk                => clk,
    reset              => reset,
    txCord             => txCord,
    iRgb               => re_05_space,
    oRgb               => re_06_space);
    
process (clk) begin
    if rising_edge(clk) then
        re_07_space <=re_06_space;
    end if;
end process;
    

    
    oRgb.red      <=re_06_space.red;
    oRgb.green    <=re_06_space.green;
    oRgb.blue     <=re_06_space.blue;
    oRgb.valid    <=re_06_space.valid;

--rgb_contrast_brightness_3_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.40,16,-3),
--    exposer_val  => 10)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_06_space,
--    oRgb              => re_07_space);
--rgb_range_3_inst: rgb_range
--generic map (
--    i_data_width       => i_data_width)
--port map (                  
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_07_space,
--    oRgb               => re_08_space);
--recolor_space_5_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_08_space,
--    oRgb               => re_09_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_6_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_09_space,
--    oRgb               => re_10_space);
--rgb_contrast_brightness_4_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(0.95,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_10_space,
--    oRgb              => re_11_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_7_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_11_space,
--    oRgb               => re_12_space);
--rgb_contrast_brightness_5_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.00,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_12_space,
--    oRgb              => re_13_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_8_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_13_space,
--    oRgb               => re_14_space);
--rgb_contrast_brightness_6_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.05,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_14_space,
--    oRgb              => re_15_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_9_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_15_space,
--    oRgb               => re_16_space);
--rgb_contrast_brightness_7_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.10,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_16_space,
--    oRgb              => re_17_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_10_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_17_space,
--    oRgb               => re_18_space);
--rgb_contrast_brightness_8_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.20,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_18_space,
--    oRgb              => re_19_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_11_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_19_space,
--    oRgb               => re_20_space);
--rgb_contrast_brightness_9_inst: rgb_contrast_brightness_level_1
--generic map (
--    contrast_val  => to_sfixed(1.30,16,-3),
--    exposer_val  => 0)
--port map (                  
--    clk               => clk,
--    rst_l             => reset,
--    iRgb              => re_20_space,
--    oRgb              => re_21_space);
--rgb_range_9_inst: rgb_range
--generic map (
--    i_data_width       => i_data_width)
--port map (                  
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_21_space,
--    oRgb               => re_22_space);
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--recolor_space_12_inst: pixel_localization
--generic map(
--    neighboring_pixel_threshold => neighboring_pixel_threshold,
--    img_width         => img_width,
--    i_data_width      => i_data_width)
--port map(
--    clk                => clk,
--    reset              => reset,
--    iRgb               => re_22_space,
--    oRgb               => re_23_space);

------------------------------------------------------------------------------
------------------------------------------------------------------------------
end behavioral;